//----------------------------------------------------------------------------
// Example
//----------------------------------------------------------------------------

module mux_4_1_width_2
(
  input  [1:0] d0, d1, d2, d3,
  input  [1:0] sel,
  output [1:0] y
);

  assign y = sel [1] ? (sel [0] ? d3 : d2)
                     : (sel [0] ? d1 : d0);

endmodule

//----------------------------------------------------------------------------
// Task
//----------------------------------------------------------------------------

module mux_4_1
(
  input  [3:0] d0, d1, d2, d3,
  input  [1:0] sel,
  output [3:0] y
);

mux_4_1_width_2 gate_1(
.d0(d0[0:1]), .d1(d1[0:1]), .d2(d2[0:1]), .d3(d3[0:1]), .sel(sel), .y(y[0:1])
);
mux_4_1_width_2 gate_2(
.d0(d0[2:3]), .d1(d1[2:3]), .d2(d2[2:3]), .d3(d3[2:3]), .sel(sel), .y(y[2:3])
);
  // Task:
  // Implement mux_4_1 with 4-bit data
  // using two instances of mux_4_1_width_2 with 2-bit data


endmodule
